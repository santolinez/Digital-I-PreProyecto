module borrar
endmodule