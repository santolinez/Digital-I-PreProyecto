//`include "Maq_Est_Y_Modos.v"

module Maq_Est_Y_Modos_TB();
    
    reg clk;
    reg reset;

    reg Boton_Comida;
    reg Boton_Medicina;

    wire sseg;
    wire an;


  
    Maq_Est_Y_Modos  uut(
        .clk(clk),
        .reset(reset),
        .Boton_Comida(Boton_Comida),
        .Boton_Medicina(Bot_Medicina)
    );

    initial begin
        clk = 0;
        reset = 0;
        Boton_Comida = 0;
        Boton_Medicina = 0;
    end 

    always #1 clk = ~clk;
    always #500 reset = ~reset;
    always #15 Boton_Comida = ~Boton_Comida;
    always #35 Boton_Medicina = ~Boton_Medicina;
  

endmodule
