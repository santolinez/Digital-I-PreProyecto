//`include "ili9341_controller.v"
//`include "freq_divider.v"


module ili9341_top #(parameter RESOLUTION = 240*240, parameter PIXEL_SIZE = 16)(
        input wire clk, //125MHz
        input wire rst,
        output wire spi_mosi,
        output wire spi_cs,
        output wire spi_sck,
        output wire spi_dc
    );

    wire clk_out;
    wire clk_input_data;
	 reg [PIXEL_SIZE-1:0] AMARILLO;
    reg [PIXEL_SIZE-1:0] current_pixel;
    reg [PIXEL_SIZE-1:0] pixel_data_mem[0:RESOLUTION/9-1];

    reg [$clog2(RESOLUTION)-1:0] pixel_counter;
	reg [1:0]counter_horizontal,counter_vertical;
    reg transmission_done;

    initial begin
        current_pixel <= 'b0;
        $readmemh("C:/Users/otro/Documents/Mecatronica/6-Sexto-Semestre/DigitalI/Proyecto/ILI/PolloBorroso_80x80.txt", pixel_data_mem);
        pixel_counter <= 'b0;
        transmission_done <= 'b0; 
        counter_horizontal <= 'b0; 
        counter_vertical <= 'b0;
    end

    freq_divider #(2) freq_divider20MHz (
        .clk(clk),
        .rst(rst),
        .clk_out(clk_out)
    );  

    always @(posedge clk_input_data) begin
        if (!rst) begin
			AMARILLO='h07FF;
            pixel_counter <= 'b0;
            current_pixel <= 'b0;
            transmission_done <= 'b0;
            counter_horizontal <= 'b0; 
            counter_vertical <= 'b0; 
        end else if (!transmission_done) begin
            if (counter_horizontal==1 )begin
                    pixel_counterM<=pixel_counterM+'b1;
            end
			if(pixel_counter==240)begin 
                counter_vertical<=counter_vertical+1;
                 if(counter_vertical==1)begin 
                pixel_counterM<=pixel_counterM+'b1;
                 end else begin
                pixel_counterM<=pixel_counterM-'d80;    
                 end
            end
                pixel_counter <= pixel_counter + 'b1;
                current_pixel <=pixel_data_mem[pixel_counterM]; //AMARILLO;
            if (pixel_counter == RESOLUTION-1) begin
                transmission_done <= 'b1; 
            end
        end
    end

    ili9341_controller ili9341(
		.clk(clk_out), 
		.rst(rst),
        .frame_done(transmission_done), 
        .input_data(current_pixel),
        .spi_mosi(spi_mosi),
		.spi_sck(spi_sck), 
        .spi_cs(spi_cs), 
        .spi_dc(spi_dc),
        .data_clk(clk_input_data)
    );

endmodule
